module bor(
    input a,
    input b,
    output r
);

    
    assign  r =a|b;
    
endmodule